library ieee;
use ieee.std_logic_1164.all;
package mem_package is
type arr is array (525 downto 0) of std_logic_vector(7 downto 0);
constant MEM_INIT : arr:= (
0 => "00000010",
1 => "00110010",
2 => "00000010",
3 => "00110100",
4 => "00000010",
5 => "00111010",
6 => "00000010",
7 => "00110110",
8 => "10000001",
9 => "01000000",
10 => "00100000",
11 => "00000000",
12 => "01000010",
13 => "01001001",
14 => "10000011",
15 => "01000000",
16 => "00110001",
17 => "00001001",
18 => "00011001",
19 => "00000010",
20 => "00010010",
21 => "00000010",
22 => "11000010",
23 => "01010000",
24 => "11000010",
25 => "01000100",
26 => "10000001",
27 => "01010110",
28 => "00000000",
29 => "10000100",
30 => "00011001",
31 => "00011110",
32 => "11011001",
33 => "00011111",
34 => "10000000",
35 => "01001001",
36 => "10100001",
37 => "00100111",
38 => "10001000",
39 => "00101011",
512 => "00000000",
513 => "00000000",
514 => "00000010",
515 => "00000000",
516 => "00000110",
517 => "00000000",
518 => "00000000",
519 => "00000001",
520 => "00000101",
521 => "00000000",
522 => "00000110",
523 => "00000000",
524 => "00000000",
525 => "00000001",
others => (others => '0'));
end package mem_package;
