library ieee;
use ieee.std_logic_1164.all;
package mem_package is
type arr is array (65535 downto 0) of std_logic_vector(7 downto 0);
constant MEM_INIT : arr:= (
0 => "00000001",
1 => "00110010",
2 => "00000001",
3 => "00110100",
4 => "00000010",
5 => "00110110",
6 => "10100000",
7 => "00000110",
8 => "11101000",
9 => "00001000",
10 => "01110000",
11 => "00101011",
12 => "01110000",
13 => "00101101",
14 => "10010001",
15 => "00000100",
16 => "10001000",
17 => "00101101",
18 => "11011001",
19 => "00000110",
20 => "00010101",
21 => "00110000",
22 => "01010000",
23 => "00000000",
24 => "10000101",
25 => "11000000",
26 => "11001000",
27 => "00100100",
28 => "10010000",
29 => "00100100",
30 => "00000010",
31 => "00110010",
32 => "00000000",
33 => "10000000",
34 => "00000000",
35 => "00110000",
36 => "00000010",
37 => "00010000",
38 => "00001010",
39 => "01011101",
40 => "00001010",
41 => "01000101",
42 => "10101000",
43 => "00000100",
44 => "01011010",
45 => "00000001",
46 => "11001101",
47 => "00010110",
48 => "00001111",
49 => "01110000",
50 => "11110000",
51 => "01100000",
52 => "00000000",
53 => "10000000",
others => (others => '0'));
end package mem_package;
